library verilog;
use verilog.vl_types.all;
entity check_d_tb is
end check_d_tb;
